`include "../basics/instruction_memory.v"

module controller ();

endmodule