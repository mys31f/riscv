`include "instruction_memory.v"

module register (
    input a1, a2, a3, wd,
    output b
);

endmodule
