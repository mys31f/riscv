module register (
    input a,
    output b
);

endmodule