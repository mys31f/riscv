module sign_extender (
    input [11:0] in_se,
    output reg [31:0] out_se
);
    
endmodule
