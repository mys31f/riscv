`include "program_counter.v"
`include "adder.v"

module instruction_memory (
    input a;
    output rd;
) 
    

endmodule