`include "./basics/adder.v"
`include "./basics/program_counter.v"
`include "./basics/instruction_memory.v"
`include "./basics/register.v"
`include "./basics/data_memory.v"
`include "./part2/controller.v"
`include "./part2/alu.v"
`include "./part2/sign_extender.v"

module cpu (
    input clk,
    input rst
)

endmodule