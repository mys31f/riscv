module data_memory (
    input [31:0] a,
    input [31:0] wd,
    input clk,
    input we,
    output [31:0] rd
);


endmodule
